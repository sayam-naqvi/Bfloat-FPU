##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Fri Jul  8 20:12:22 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_proj_example
  CLASS BLOCK ;
  SIZE 818.340000 BY 814.640000 ;
  FOREIGN user_proj_example 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5831 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 152.038 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 811.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.852 LAYER met3  ;
    ANTENNAMAXAREACAR 179.059 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 954.839 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.107277 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1.605000 0.000000 1.745000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 90.006 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.611 LAYER met2  ;
    ANTENNAMAXAREACAR 13.992 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.6911 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.620000 0.000000 0.760000 0.490000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.920000 0.000000 174.060000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.485000 0.000000 58.625000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.595000 0.000000 175.735000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.250000 0.000000 172.390000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.575000 0.000000 170.715000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.905000 0.000000 169.045000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.230000 0.000000 167.370000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.020000 0.000000 112.160000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.350000 0.000000 110.490000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.675000 0.000000 108.815000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.000000 0.000000 107.140000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.330000 0.000000 105.470000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.655000 0.000000 103.795000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.985000 0.000000 102.125000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.310000 0.000000 100.450000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.635000 0.000000 98.775000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.965000 0.000000 97.105000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.290000 0.000000 95.430000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.620000 0.000000 93.760000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.945000 0.000000 92.085000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.270000 0.000000 90.410000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.600000 0.000000 88.740000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.925000 0.000000 87.065000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.255000 0.000000 85.395000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.580000 0.000000 83.720000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.905000 0.000000 82.045000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.235000 0.000000 80.375000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.560000 0.000000 78.700000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.890000 0.000000 77.030000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.215000 0.000000 75.355000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.540000 0.000000 73.680000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.870000 0.000000 72.010000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.195000 0.000000 70.335000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.525000 0.000000 68.665000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.850000 0.000000 66.990000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.175000 0.000000 65.315000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.505000 0.000000 63.645000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.830000 0.000000 61.970000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.160000 0.000000 60.300000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.810000 0.000000 56.950000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.140000 0.000000 55.280000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.465000 0.000000 53.605000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.795000 0.000000 51.935000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.120000 0.000000 50.260000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.445000 0.000000 48.585000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.775000 0.000000 46.915000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.100000 0.000000 45.240000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.430000 0.000000 43.570000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.755000 0.000000 41.895000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.080000 0.000000 40.220000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.410000 0.000000 38.550000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.735000 0.000000 36.875000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.065000 0.000000 35.205000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.390000 0.000000 33.530000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.715000 0.000000 31.855000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.045000 0.000000 30.185000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.370000 0.000000 28.510000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.700000 0.000000 26.840000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.025000 0.000000 25.165000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.350000 0.000000 23.490000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.680000 0.000000 21.820000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.005000 0.000000 20.145000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.335000 0.000000 18.475000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.660000 0.000000 16.800000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.985000 0.000000 15.125000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.315000 0.000000 13.455000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.640000 0.000000 11.780000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.970000 0.000000 10.110000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.295000 0.000000 8.435000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.620000 0.000000 6.760000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.950000 0.000000 5.090000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 3.275000 0.000000 3.415000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 165.555000 0.000000 165.695000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 163.885000 0.000000 164.025000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 358.3 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7944 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.837 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 162.210000 0.000000 162.350000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 160.540000 0.000000 160.680000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 158.865000 0.000000 159.005000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 157.190000 0.000000 157.330000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 155.520000 0.000000 155.660000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 153.845000 0.000000 153.985000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 152.175000 0.000000 152.315000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 150.500000 0.000000 150.640000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 148.825000 0.000000 148.965000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 147.155000 0.000000 147.295000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 145.480000 0.000000 145.620000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 358.3 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7944 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.837 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 143.810000 0.000000 143.950000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 142.135000 0.000000 142.275000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 358.3 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7944 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.837 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 140.460000 0.000000 140.600000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 138.790000 0.000000 138.930000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 137.115000 0.000000 137.255000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 135.445000 0.000000 135.585000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 133.770000 0.000000 133.910000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 132.095000 0.000000 132.235000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 130.425000 0.000000 130.565000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 128.750000 0.000000 128.890000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 127.080000 0.000000 127.220000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 125.405000 0.000000 125.545000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 123.730000 0.000000 123.870000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 358.3 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7944 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.837 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 122.060000 0.000000 122.200000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 358.033 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7944 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.57 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 120.385000 0.000000 120.525000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 358.033 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7944 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.57 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 118.715000 0.000000 118.855000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 358.033 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7944 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.57 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 117.040000 0.000000 117.180000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 358.033 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7944 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.57 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 115.365000 0.000000 115.505000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 75.2061 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 364.623 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.89008 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 96.6168 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 498.16 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.89008 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 113.695000 0.000000 113.835000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.740000 0.000000 389.880000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.065000 0.000000 388.205000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.395000 0.000000 386.535000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.720000 0.000000 384.860000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.045000 0.000000 383.185000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.375000 0.000000 381.515000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.700000 0.000000 379.840000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.030000 0.000000 378.170000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.355000 0.000000 376.495000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.680000 0.000000 374.820000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.010000 0.000000 373.150000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.335000 0.000000 371.475000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.665000 0.000000 369.805000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.990000 0.000000 368.130000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.315000 0.000000 366.455000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.645000 0.000000 364.785000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.970000 0.000000 363.110000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.300000 0.000000 361.440000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.625000 0.000000 359.765000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.950000 0.000000 358.090000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.280000 0.000000 356.420000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.605000 0.000000 354.745000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.935000 0.000000 353.075000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.260000 0.000000 351.400000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.585000 0.000000 349.725000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.915000 0.000000 348.055000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.240000 0.000000 346.380000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.570000 0.000000 344.710000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.895000 0.000000 343.035000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.220000 0.000000 341.360000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.550000 0.000000 339.690000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.875000 0.000000 338.015000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.205000 0.000000 336.345000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.530000 0.000000 334.670000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.855000 0.000000 332.995000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.185000 0.000000 331.325000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.510000 0.000000 329.650000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.840000 0.000000 327.980000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.165000 0.000000 326.305000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.490000 0.000000 324.630000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.820000 0.000000 322.960000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.145000 0.000000 321.285000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.475000 0.000000 319.615000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.800000 0.000000 317.940000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.125000 0.000000 316.265000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.455000 0.000000 314.595000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.780000 0.000000 312.920000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.110000 0.000000 311.250000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.435000 0.000000 309.575000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.760000 0.000000 307.900000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.090000 0.000000 306.230000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.415000 0.000000 304.555000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.745000 0.000000 302.885000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.070000 0.000000 301.210000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.395000 0.000000 299.535000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.725000 0.000000 297.865000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.050000 0.000000 296.190000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.380000 0.000000 294.520000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.705000 0.000000 292.845000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.030000 0.000000 291.170000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.360000 0.000000 289.500000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.685000 0.000000 287.825000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.9456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.567 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 64.5333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 345.584 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 19.305 LAYER met3  ;
    ANTENNAMAXAREACAR 5.86818 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 28.6094 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0960331 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 286.015000 0.000000 286.155000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.8145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 219.881 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1180.21 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 10.62 LAYER met4  ;
    ANTENNAMAXAREACAR 108.334 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 543.766 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 284.340000 0.000000 284.480000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.665000 0.000000 282.805000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.995000 0.000000 281.135000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.320000 0.000000 279.460000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.650000 0.000000 277.790000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.975000 0.000000 276.115000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.300000 0.000000 274.440000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.630000 0.000000 272.770000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.955000 0.000000 271.095000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.285000 0.000000 269.425000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.610000 0.000000 267.750000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.935000 0.000000 266.075000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.265000 0.000000 264.405000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.590000 0.000000 262.730000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.920000 0.000000 261.060000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.245000 0.000000 259.385000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.570000 0.000000 257.710000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.900000 0.000000 256.040000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.225000 0.000000 254.365000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.555000 0.000000 252.695000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.880000 0.000000 251.020000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.205000 0.000000 249.345000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.535000 0.000000 247.675000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.860000 0.000000 246.000000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.190000 0.000000 244.330000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.515000 0.000000 242.655000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.840000 0.000000 240.980000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.170000 0.000000 239.310000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.495000 0.000000 237.635000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.825000 0.000000 235.965000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.150000 0.000000 234.290000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.475000 0.000000 232.615000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.805000 0.000000 230.945000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.809 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.937 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8052 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.1905 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.318651 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.130000 0.000000 229.270000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.83 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 21.482 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.9551 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 227.460000 0.000000 227.600000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2515 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 27.1295 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 122.241 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 225.785000 0.000000 225.925000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2124 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.836 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 11.7596 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.1798 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 224.110000 0.000000 224.250000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1438 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.493 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 9.71434 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.7273 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 222.440000 0.000000 222.580000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.7415 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.813 LAYER met2  ;
    ANTENNAMAXAREACAR 6.78874 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.6122 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 220.765000 0.000000 220.905000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3388 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.478 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 10.8687 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 48.4909 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 219.095000 0.000000 219.235000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6792 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 8.40509 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.132 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.289606 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 217.420000 0.000000 217.560000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1775 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6715 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 5.47576 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.2172 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 215.745000 0.000000 215.885000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0503 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0255 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 9.46404 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.4758 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 214.075000 0.000000 214.215000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5108 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.22 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.08997 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.7758 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 212.400000 0.000000 212.540000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.59 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.724 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 11.9871 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.4465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 210.730000 0.000000 210.870000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 18.2282 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.2682 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.055000 0.000000 209.195000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.826 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.74397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.8963 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.147071 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 207.380000 0.000000 207.520000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0912 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.122 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 6.30707 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.6889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 205.710000 0.000000 205.850000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8764 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.221 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.7748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.57239 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.8889 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.352458 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 204.035000 0.000000 204.175000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.365000 0.000000 202.505000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.690000 0.000000 200.830000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.015000 0.000000 199.155000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.345000 0.000000 197.485000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.670000 0.000000 195.810000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.000000 0.000000 194.140000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.325000 0.000000 192.465000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.650000 0.000000 190.790000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.980000 0.000000 189.120000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.305000 0.000000 187.445000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.635000 0.000000 185.775000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.960000 0.000000 184.100000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.285000 0.000000 182.425000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.615000 0.000000 180.755000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4372 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.96 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 55.7155 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 276.281 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 178.940000 0.000000 179.080000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.270000 0.000000 177.410000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3509 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.3045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 603.885000 0.000000 604.025000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.406 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 602.210000 0.000000 602.350000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.406 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 600.535000 0.000000 600.675000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.3535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 598.865000 0.000000 599.005000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.406 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 597.190000 0.000000 597.330000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.406 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 595.520000 0.000000 595.660000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.3535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 593.845000 0.000000 593.985000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.406 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 592.170000 0.000000 592.310000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.3535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 590.500000 0.000000 590.640000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.3535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 588.825000 0.000000 588.965000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.3535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 587.155000 0.000000 587.295000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.406 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 585.480000 0.000000 585.620000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.3535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 583.805000 0.000000 583.945000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.3535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 582.135000 0.000000 582.275000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.406 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 580.460000 0.000000 580.600000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3901 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.5775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 578.790000 0.000000 578.930000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3509 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.3045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.6383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 577.115000 0.000000 577.255000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1734 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.631 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.49 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 575.440000 0.000000 575.580000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 573.770000 0.000000 573.910000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 572.095000 0.000000 572.235000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 570.425000 0.000000 570.565000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 568.750000 0.000000 568.890000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 567.075000 0.000000 567.215000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 565.405000 0.000000 565.545000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 563.730000 0.000000 563.870000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 562.060000 0.000000 562.200000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 560.385000 0.000000 560.525000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 558.710000 0.000000 558.850000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 557.040000 0.000000 557.180000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 555.365000 0.000000 555.505000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 553.695000 0.000000 553.835000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 552.020000 0.000000 552.160000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 550.345000 0.000000 550.485000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 548.675000 0.000000 548.815000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 547.000000 0.000000 547.140000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 545.330000 0.000000 545.470000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 543.655000 0.000000 543.795000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 541.980000 0.000000 542.120000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 540.310000 0.000000 540.450000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 538.635000 0.000000 538.775000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 536.965000 0.000000 537.105000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 535.290000 0.000000 535.430000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 533.615000 0.000000 533.755000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 531.945000 0.000000 532.085000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 530.270000 0.000000 530.410000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 528.600000 0.000000 528.740000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 526.925000 0.000000 527.065000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 525.250000 0.000000 525.390000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 523.580000 0.000000 523.720000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 521.905000 0.000000 522.045000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 520.235000 0.000000 520.375000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 518.560000 0.000000 518.700000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 516.885000 0.000000 517.025000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 515.215000 0.000000 515.355000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 513.540000 0.000000 513.680000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 511.870000 0.000000 512.010000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 510.195000 0.000000 510.335000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 508.520000 0.000000 508.660000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 506.850000 0.000000 506.990000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 505.175000 0.000000 505.315000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 503.505000 0.000000 503.645000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 501.830000 0.000000 501.970000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 500.155000 0.000000 500.295000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 498.485000 0.000000 498.625000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 496.810000 0.000000 496.950000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 495.140000 0.000000 495.280000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 493.465000 0.000000 493.605000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 491.790000 0.000000 491.930000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 490.120000 0.000000 490.260000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 488.445000 0.000000 488.585000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 486.775000 0.000000 486.915000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 485.100000 0.000000 485.240000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 483.425000 0.000000 483.565000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 481.755000 0.000000 481.895000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 480.080000 0.000000 480.220000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 478.410000 0.000000 478.550000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 476.735000 0.000000 476.875000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 475.060000 0.000000 475.200000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 473.390000 0.000000 473.530000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1734 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.631 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.49 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 471.715000 0.000000 471.855000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6141 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.9095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.191 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.431 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.5968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.32 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 470.045000 0.000000 470.185000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.617 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7155 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.6208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 190.448 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 468.370000 0.000000 468.510000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1805 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.721 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.431 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.6728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 233.392 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 466.695000 0.000000 466.835000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.371 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.93 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7155 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.7738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.264 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 465.025000 0.000000 465.165000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9022 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.35 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7155 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.4638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 210.944 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 463.350000 0.000000 463.490000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8115 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.482 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7155 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.6778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 158.752 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 461.680000 0.000000 461.820000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.2973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 96.2605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 460.005000 0.000000 460.145000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.9924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 99.736 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 458.330000 0.000000 458.470000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.341 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7155 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.8848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.856 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 456.660000 0.000000 456.800000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.25 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 161.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7155 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.3988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.264 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 454.985000 0.000000 455.125000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.6065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.8065 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 453.315000 0.000000 453.455000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6047 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 173.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.431 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.1438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 171.904 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 451.640000 0.000000 451.780000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6509 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.52 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 179.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.1438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 171.904 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 449.965000 0.000000 450.105000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.6337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.9425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 448.295000 0.000000 448.435000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.8416 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 93.982 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 446.620000 0.000000 446.760000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.4345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.313 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 178.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.4948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.776 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 444.950000 0.000000 445.090000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1734 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.631 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.49 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 443.275000 0.000000 443.415000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 441.600000 0.000000 441.740000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 439.930000 0.000000 440.070000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 438.255000 0.000000 438.395000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 436.585000 0.000000 436.725000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 434.910000 0.000000 435.050000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 433.235000 0.000000 433.375000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 431.565000 0.000000 431.705000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 429.890000 0.000000 430.030000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.1832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 113.536 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 566.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 428.220000 0.000000 428.360000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.2028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.802 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 115.18 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 570.84 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.241315 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 426.545000 0.000000 426.685000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 424.870000 0.000000 425.010000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 423.200000 0.000000 423.340000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 421.525000 0.000000 421.665000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 419.855000 0.000000 419.995000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 418.180000 0.000000 418.320000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 416.505000 0.000000 416.645000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 414.835000 0.000000 414.975000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 413.160000 0.000000 413.300000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 411.490000 0.000000 411.630000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 409.815000 0.000000 409.955000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 408.140000 0.000000 408.280000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 406.470000 0.000000 406.610000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 404.795000 0.000000 404.935000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 403.125000 0.000000 403.265000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 401.450000 0.000000 401.590000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 399.775000 0.000000 399.915000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 398.105000 0.000000 398.245000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 396.430000 0.000000 396.570000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 358.3 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7944 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.837 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 394.760000 0.000000 394.900000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 358.033 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7944 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.57 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 393.085000 0.000000 393.225000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 73.3338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.24 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 94.7445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.6285 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 391.410000 0.000000 391.550000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.660000 0.000000 816.800000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.355000 0.000000 816.495000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.680000 0.000000 814.820000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.010000 0.000000 813.150000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.335000 0.000000 811.475000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.660000 0.000000 809.800000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.990000 0.000000 808.130000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.315000 0.000000 806.455000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.645000 0.000000 804.785000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.970000 0.000000 803.110000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.295000 0.000000 801.435000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.625000 0.000000 799.765000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.950000 0.000000 798.090000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.280000 0.000000 796.420000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.605000 0.000000 794.745000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.930000 0.000000 793.070000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.260000 0.000000 791.400000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.585000 0.000000 789.725000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.915000 0.000000 788.055000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.240000 0.000000 786.380000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.565000 0.000000 784.705000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.895000 0.000000 783.035000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.220000 0.000000 781.360000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.550000 0.000000 779.690000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.875000 0.000000 778.015000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.200000 0.000000 776.340000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.530000 0.000000 774.670000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.855000 0.000000 772.995000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.185000 0.000000 771.325000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.510000 0.000000 769.650000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.835000 0.000000 767.975000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.165000 0.000000 766.305000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.490000 0.000000 764.630000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.820000 0.000000 762.960000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.145000 0.000000 761.285000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.470000 0.000000 759.610000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.800000 0.000000 757.940000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.125000 0.000000 756.265000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.455000 0.000000 754.595000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.780000 0.000000 752.920000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.105000 0.000000 751.245000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.435000 0.000000 749.575000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.760000 0.000000 747.900000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.090000 0.000000 746.230000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.415000 0.000000 744.555000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.740000 0.000000 742.880000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.070000 0.000000 741.210000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.395000 0.000000 739.535000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.725000 0.000000 737.865000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.050000 0.000000 736.190000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.375000 0.000000 734.515000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.705000 0.000000 732.845000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030000 0.000000 731.170000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.360000 0.000000 729.500000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.685000 0.000000 727.825000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.010000 0.000000 726.150000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.340000 0.000000 724.480000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.665000 0.000000 722.805000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.995000 0.000000 721.135000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.320000 0.000000 719.460000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.645000 0.000000 717.785000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.975000 0.000000 716.115000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7231 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 55.792 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 298.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.0584 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 295.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 33.966 LAYER met4  ;
    ANTENNAMAXAREACAR 6.58664 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 22.0302 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.346263 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 714.300000 0.000000 714.440000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8114 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.896 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 50.7659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 271.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.479 LAYER met3  ;
    ANTENNAMAXAREACAR 48.3481 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 249.855 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.177688 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 218.769 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1170.05 LAYER met4  ;
    ANTENNAGATEAREA 16.35 LAYER met4  ;
    ANTENNAMAXAREACAR 107.411 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 542.732 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 712.630000 0.000000 712.770000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.955000 0.000000 711.095000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.280000 0.000000 709.420000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.610000 0.000000 707.750000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.935000 0.000000 706.075000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.265000 0.000000 704.405000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.590000 0.000000 702.730000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.915000 0.000000 701.055000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.245000 0.000000 699.385000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.570000 0.000000 697.710000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.900000 0.000000 696.040000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.225000 0.000000 694.365000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.550000 0.000000 692.690000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.880000 0.000000 691.020000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.205000 0.000000 689.345000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.535000 0.000000 687.675000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.860000 0.000000 686.000000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3825 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 2.33525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.5232 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 684.185000 0.000000 684.325000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.318 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 2.57995 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.4187 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 682.515000 0.000000 682.655000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6512 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.148 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 2.11303 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.19747 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 680.840000 0.000000 680.980000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5966 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.875 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 2.45641 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.8793 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 679.170000 0.000000 679.310000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0225 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 3.00556 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.8747 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 677.495000 0.000000 677.635000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4492 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.138 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 3.18889 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.4116 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 675.820000 0.000000 675.960000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5619 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7015 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 3.20434 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.6222 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 674.150000 0.000000 674.290000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7138 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.461 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 3.36687 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.3985 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 672.475000 0.000000 672.615000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.47434 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.6808 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 670.805000 0.000000 670.945000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.821 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.59899 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.4717 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 669.130000 0.000000 669.270000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0089 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9365 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.70202 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.0283 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 667.455000 0.000000 667.595000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9837 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8105 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.97354 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.5556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 665.785000 0.000000 665.925000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.302 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 3.41495 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.9217 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 664.110000 0.000000 664.250000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.847 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 2.74773 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.1894 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 662.440000 0.000000 662.580000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0955 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 2.10242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.14444 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 660.765000 0.000000 660.905000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.239 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 2.12232 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.2803 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 659.090000 0.000000 659.230000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.568 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 24.9749 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 118.212 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 657.420000 0.000000 657.560000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9319 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5515 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.60525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.0182 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 655.745000 0.000000 655.885000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0509 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1465 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.586 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.6808 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 654.075000 0.000000 654.215000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.996 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.3358 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.0162 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 652.400000 0.000000 652.540000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9669 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7265 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.2218 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.0808 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 650.725000 0.000000 650.865000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6757 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2705 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.87111 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.3475 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 649.055000 0.000000 649.195000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4916 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.35 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.0967 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.2343 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 647.380000 0.000000 647.520000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.469 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.07434 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.7091 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 645.710000 0.000000 645.850000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4429 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.1065 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 12.4505 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.2444 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 644.035000 0.000000 644.175000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.424 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 12.6591 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.0465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 642.360000 0.000000 642.500000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2826 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.305 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 11.6537 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.6061 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 640.690000 0.000000 640.830000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6935 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 11.0893 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.6909 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 639.015000 0.000000 639.155000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.7931 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.9576 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 637.345000 0.000000 637.485000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.525 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.8094 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.798 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 635.670000 0.000000 635.810000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1165 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.2218 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.0808 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 633.995000 0.000000 634.135000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 14.1523 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.7899 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 632.325000 0.000000 632.465000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.650000 0.000000 630.790000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.980000 0.000000 629.120000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.305000 0.000000 627.445000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.630000 0.000000 625.770000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.960000 0.000000 624.100000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.285000 0.000000 622.425000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.615000 0.000000 620.755000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.940000 0.000000 619.080000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.265000 0.000000 617.405000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.595000 0.000000 615.735000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.920000 0.000000 614.060000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.250000 0.000000 612.390000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.575000 0.000000 610.715000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.900000 0.000000 609.040000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.001 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 15.7723 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.0879 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 607.230000 0.000000 607.370000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.555000 0.000000 605.695000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 39.590000 0.800000 39.890000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 99.195000 0.800000 99.495000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 158.800000 0.800000 159.100000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 218.410000 0.800000 218.710000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 278.015000 0.800000 278.315000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 337.625000 0.800000 337.925000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 397.230000 0.800000 397.530000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 456.835000 0.800000 457.135000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 516.445000 0.800000 516.745000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 576.050000 0.800000 576.350000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 635.660000 0.800000 635.960000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 695.265000 0.800000 695.565000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 754.870000 0.800000 755.170000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 810.540000 0.800000 810.840000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.880000 814.150000 63.020000 814.640000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.300000 814.150000 157.440000 814.640000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.720000 814.150000 251.860000 814.640000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.145000 814.150000 346.285000 814.640000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.565000 814.150000 440.705000 814.640000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.990000 814.150000 535.130000 814.640000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.410000 814.150000 629.550000 814.640000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.830000 814.150000 723.970000 814.640000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.680000 814.150000 810.820000 814.640000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 777.440000 818.340000 777.740000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 721.895000 818.340000 722.195000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 666.355000 818.340000 666.655000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 610.810000 818.340000 611.110000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 555.270000 818.340000 555.570000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 499.730000 818.340000 500.030000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 444.185000 818.340000 444.485000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 388.645000 818.340000 388.945000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 333.100000 818.340000 333.400000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 57.7414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 308.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 15.1168 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 80.0687 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 277.560000 818.340000 277.860000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 222.020000 818.340000 222.320000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 166.475000 818.340000 166.775000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 110.935000 818.340000 111.235000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 55.390000 818.340000 55.690000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.540000 9.610000 818.340000 9.910000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 20.8 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 130.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 19.720000 0.800000 20.020000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0122 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 20.4183 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 128.244 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 79.325000 0.800000 79.625000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0122 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 20.4183 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 128.244 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 138.935000 0.800000 139.235000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0122 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 20.4183 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 128.244 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 198.540000 0.800000 198.840000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 258.145000 0.800000 258.445000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 317.755000 0.800000 318.055000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 377.360000 0.800000 377.660000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.9446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.5521 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.117 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 436.970000 0.800000 437.270000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 496.575000 0.800000 496.875000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 556.180000 0.800000 556.480000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 615.790000 0.800000 616.090000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 675.395000 0.800000 675.695000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 735.005000 0.800000 735.305000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 794.610000 0.800000 794.910000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3406 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 81.424 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 70.9068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 378.64 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 31.405000 814.150000 31.545000 814.640000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.375 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.596 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 2.862 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 61.4808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 328.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 125.825000 814.150000 125.965000 814.640000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3141 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.154 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 74.4018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 397.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 220.250000 814.150000 220.390000 814.640000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 159.115 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 849.552 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 314.670000 814.150000 314.810000 814.640000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.3858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.736 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 2.673 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 174.784 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 266.016 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 409.090000 814.150000 409.230000 814.640000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.2162 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 235.802 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.57 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 65.1798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 348.096 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 503.515000 814.150000 503.655000 814.640000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.875 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.214 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.431 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 135.898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 725.728 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 597.935000 814.150000 598.075000 814.640000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4467 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.0725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 145.001 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 773.808 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 692.360000 814.150000 692.500000 814.640000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.5705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 72.6915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 46.147 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 246.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 142.16 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 758.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 786.780000 814.150000 786.920000 814.640000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 40.0486 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 213.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.862 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 172.681 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 921.904 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 795.950000 818.340000 796.250000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.1606 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 208.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 158.087 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 844.544 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 740.410000 818.340000 740.710000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 141.007 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 752.976 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 684.870000 818.340000 685.170000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9471 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 127.933 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 683.248 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 629.325000 818.340000 629.625000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5611 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 116.779 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 623.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 573.785000 818.340000 574.085000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.7414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 260.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.4346 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 216.592 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 518.240000 818.340000 518.540000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.3064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 194.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.431 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.9168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 277.36 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 462.700000 818.340000 463.000000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 407.160000 818.340000 407.460000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.623 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 351.615000 818.340000 351.915000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8271 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 296.075000 818.340000 296.375000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5466 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 240.530000 818.340000 240.830000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 184.990000 818.340000 185.290000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4433 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 129.450000 818.340000 129.750000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.5183 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 73.905000 818.340000 74.205000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4433 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 18.365000 818.340000 18.665000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 20.8 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 130.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 10.220000 0.800000 10.520000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 20.8 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 130.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 59.455000 0.800000 59.755000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0122 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 20.4183 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 128.244 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 119.065000 0.800000 119.365000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0122 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 20.4183 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 128.244 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 178.670000 0.800000 178.970000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.9446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.5521 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.117 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 238.280000 0.800000 238.580000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 297.885000 0.800000 298.185000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 357.490000 0.800000 357.790000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.9446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.5521 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.117 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 417.100000 0.800000 417.400000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.9446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.5521 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.117 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 476.705000 0.800000 477.005000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 536.315000 0.800000 536.615000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 595.920000 0.800000 596.220000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 655.525000 0.800000 655.825000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 715.135000 0.800000 715.435000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 774.740000 0.800000 775.040000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.0503 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.893 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.92 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 80.1155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 494.122 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 10.280000 814.150000 10.420000 814.640000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.0566 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.924 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.92 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 80.1155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 494.122 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 94.350000 814.150000 94.490000 814.640000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.0321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.802 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.92 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 80.1155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 494.122 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 188.775000 814.150000 188.915000 814.640000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.0566 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.924 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.92 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 80.1155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 494.122 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 283.195000 814.150000 283.335000 814.640000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.0321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.802 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.92 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 80.1155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 494.122 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 377.620000 814.150000 377.760000 814.640000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.0321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.802 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.92 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 80.1155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 494.122 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 472.040000 814.150000 472.180000 814.640000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.0321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.802 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.92 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 80.1155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 494.122 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 566.460000 814.150000 566.600000 814.640000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.0566 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.924 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.92 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 80.1155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 494.122 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 660.885000 814.150000 661.025000 814.640000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.0223 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.92 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 80.1155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 494.122 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 755.305000 814.150000 755.445000 814.640000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.9446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.5521 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.117 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 809.930000 818.340000 810.230000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.9446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.5521 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.117 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 758.925000 818.340000 759.225000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 703.380000 818.340000 703.680000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.9446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 109.127 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 632.296 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.804695 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 647.840000 818.340000 648.140000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8246 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 78.9887 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 485.859 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 592.300000 818.340000 592.600000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.239 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 536.755000 818.340000 537.055000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4881 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 481.215000 818.340000 481.515000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 425.670000 818.340000 425.970000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.713 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 370.130000 818.340000 370.430000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.7316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 80.6644 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 434.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.544 LAYER met4  ;
    ANTENNAMAXAREACAR 87.7046 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 462.043 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.0869 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 314.590000 818.340000 314.890000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6321 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 259.045000 818.340000 259.345000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.689 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 203.505000 818.340000 203.805000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4433 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 147.960000 818.340000 148.260000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.5183 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 92.420000 818.340000 92.720000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4433 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4509 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 817.540000 36.880000 818.340000 37.180000 ;
    END
  END io_oeb[0]
  PIN irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.0552 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.941 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.92 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 80.1155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 494.122 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1.080000 814.155000 1.220000 814.640000 ;
    END
  END irq[2]
  PIN irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.0426 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.854 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.92 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 80.1155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 494.122 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.620000 814.155000 0.760000 814.640000 ;
    END
  END irq[1]
  PIN irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.0552 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.941 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.92 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 80.1155 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 494.122 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.160000 814.155000 0.300000 814.640000 ;
    END
  END irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.560000 0.600000 2.560000 814.040000 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.780000 0.600000 817.780000 814.040000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 502.060000 388.790000 503.800000 783.570000 ;
      LAYER met4 ;
        RECT 26.740000 388.790000 28.480000 783.570000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 7.560000 7.600000 9.560000 807.040000 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.780000 7.600000 810.780000 807.040000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 30.140000 392.190000 31.880000 780.170000 ;
      LAYER met4 ;
        RECT 498.660000 392.190000 500.400000 780.170000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 818.340000 814.640000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 818.340000 814.640000 ;
    LAYER met2 ;
      RECT 1.360000 814.015000 10.140000 814.640000 ;
      RECT 0.900000 814.015000 0.940000 814.640000 ;
      RECT 0.440000 814.015000 0.480000 814.640000 ;
      RECT 0.000000 814.015000 0.020000 814.640000 ;
      RECT 810.960000 814.010000 818.340000 814.640000 ;
      RECT 787.060000 814.010000 810.540000 814.640000 ;
      RECT 755.585000 814.010000 786.640000 814.640000 ;
      RECT 724.110000 814.010000 755.165000 814.640000 ;
      RECT 692.640000 814.010000 723.690000 814.640000 ;
      RECT 661.165000 814.010000 692.220000 814.640000 ;
      RECT 629.690000 814.010000 660.745000 814.640000 ;
      RECT 598.215000 814.010000 629.270000 814.640000 ;
      RECT 566.740000 814.010000 597.795000 814.640000 ;
      RECT 535.270000 814.010000 566.320000 814.640000 ;
      RECT 503.795000 814.010000 534.850000 814.640000 ;
      RECT 472.320000 814.010000 503.375000 814.640000 ;
      RECT 440.845000 814.010000 471.900000 814.640000 ;
      RECT 409.370000 814.010000 440.425000 814.640000 ;
      RECT 377.900000 814.010000 408.950000 814.640000 ;
      RECT 346.425000 814.010000 377.480000 814.640000 ;
      RECT 314.950000 814.010000 346.005000 814.640000 ;
      RECT 283.475000 814.010000 314.530000 814.640000 ;
      RECT 252.000000 814.010000 283.055000 814.640000 ;
      RECT 220.530000 814.010000 251.580000 814.640000 ;
      RECT 189.055000 814.010000 220.110000 814.640000 ;
      RECT 157.580000 814.010000 188.635000 814.640000 ;
      RECT 126.105000 814.010000 157.160000 814.640000 ;
      RECT 94.630000 814.010000 125.685000 814.640000 ;
      RECT 63.160000 814.010000 94.210000 814.640000 ;
      RECT 31.685000 814.010000 62.740000 814.640000 ;
      RECT 10.560000 814.010000 31.265000 814.640000 ;
      RECT 0.000000 814.010000 10.140000 814.015000 ;
      RECT 0.000000 0.630000 818.340000 814.010000 ;
      RECT 816.940000 0.000000 818.340000 0.630000 ;
      RECT 814.960000 0.000000 816.215000 0.630000 ;
      RECT 813.290000 0.000000 814.540000 0.630000 ;
      RECT 811.615000 0.000000 812.870000 0.630000 ;
      RECT 809.940000 0.000000 811.195000 0.630000 ;
      RECT 808.270000 0.000000 809.520000 0.630000 ;
      RECT 806.595000 0.000000 807.850000 0.630000 ;
      RECT 804.925000 0.000000 806.175000 0.630000 ;
      RECT 803.250000 0.000000 804.505000 0.630000 ;
      RECT 801.575000 0.000000 802.830000 0.630000 ;
      RECT 799.905000 0.000000 801.155000 0.630000 ;
      RECT 798.230000 0.000000 799.485000 0.630000 ;
      RECT 796.560000 0.000000 797.810000 0.630000 ;
      RECT 794.885000 0.000000 796.140000 0.630000 ;
      RECT 793.210000 0.000000 794.465000 0.630000 ;
      RECT 791.540000 0.000000 792.790000 0.630000 ;
      RECT 789.865000 0.000000 791.120000 0.630000 ;
      RECT 788.195000 0.000000 789.445000 0.630000 ;
      RECT 786.520000 0.000000 787.775000 0.630000 ;
      RECT 784.845000 0.000000 786.100000 0.630000 ;
      RECT 783.175000 0.000000 784.425000 0.630000 ;
      RECT 781.500000 0.000000 782.755000 0.630000 ;
      RECT 779.830000 0.000000 781.080000 0.630000 ;
      RECT 778.155000 0.000000 779.410000 0.630000 ;
      RECT 776.480000 0.000000 777.735000 0.630000 ;
      RECT 774.810000 0.000000 776.060000 0.630000 ;
      RECT 773.135000 0.000000 774.390000 0.630000 ;
      RECT 771.465000 0.000000 772.715000 0.630000 ;
      RECT 769.790000 0.000000 771.045000 0.630000 ;
      RECT 768.115000 0.000000 769.370000 0.630000 ;
      RECT 766.445000 0.000000 767.695000 0.630000 ;
      RECT 764.770000 0.000000 766.025000 0.630000 ;
      RECT 763.100000 0.000000 764.350000 0.630000 ;
      RECT 761.425000 0.000000 762.680000 0.630000 ;
      RECT 759.750000 0.000000 761.005000 0.630000 ;
      RECT 758.080000 0.000000 759.330000 0.630000 ;
      RECT 756.405000 0.000000 757.660000 0.630000 ;
      RECT 754.735000 0.000000 755.985000 0.630000 ;
      RECT 753.060000 0.000000 754.315000 0.630000 ;
      RECT 751.385000 0.000000 752.640000 0.630000 ;
      RECT 749.715000 0.000000 750.965000 0.630000 ;
      RECT 748.040000 0.000000 749.295000 0.630000 ;
      RECT 746.370000 0.000000 747.620000 0.630000 ;
      RECT 744.695000 0.000000 745.950000 0.630000 ;
      RECT 743.020000 0.000000 744.275000 0.630000 ;
      RECT 741.350000 0.000000 742.600000 0.630000 ;
      RECT 739.675000 0.000000 740.930000 0.630000 ;
      RECT 738.005000 0.000000 739.255000 0.630000 ;
      RECT 736.330000 0.000000 737.585000 0.630000 ;
      RECT 734.655000 0.000000 735.910000 0.630000 ;
      RECT 732.985000 0.000000 734.235000 0.630000 ;
      RECT 731.310000 0.000000 732.565000 0.630000 ;
      RECT 729.640000 0.000000 730.890000 0.630000 ;
      RECT 727.965000 0.000000 729.220000 0.630000 ;
      RECT 726.290000 0.000000 727.545000 0.630000 ;
      RECT 724.620000 0.000000 725.870000 0.630000 ;
      RECT 722.945000 0.000000 724.200000 0.630000 ;
      RECT 721.275000 0.000000 722.525000 0.630000 ;
      RECT 719.600000 0.000000 720.855000 0.630000 ;
      RECT 717.925000 0.000000 719.180000 0.630000 ;
      RECT 716.255000 0.000000 717.505000 0.630000 ;
      RECT 714.580000 0.000000 715.835000 0.630000 ;
      RECT 712.910000 0.000000 714.160000 0.630000 ;
      RECT 711.235000 0.000000 712.490000 0.630000 ;
      RECT 709.560000 0.000000 710.815000 0.630000 ;
      RECT 707.890000 0.000000 709.140000 0.630000 ;
      RECT 706.215000 0.000000 707.470000 0.630000 ;
      RECT 704.545000 0.000000 705.795000 0.630000 ;
      RECT 702.870000 0.000000 704.125000 0.630000 ;
      RECT 701.195000 0.000000 702.450000 0.630000 ;
      RECT 699.525000 0.000000 700.775000 0.630000 ;
      RECT 697.850000 0.000000 699.105000 0.630000 ;
      RECT 696.180000 0.000000 697.430000 0.630000 ;
      RECT 694.505000 0.000000 695.760000 0.630000 ;
      RECT 692.830000 0.000000 694.085000 0.630000 ;
      RECT 691.160000 0.000000 692.410000 0.630000 ;
      RECT 689.485000 0.000000 690.740000 0.630000 ;
      RECT 687.815000 0.000000 689.065000 0.630000 ;
      RECT 686.140000 0.000000 687.395000 0.630000 ;
      RECT 684.465000 0.000000 685.720000 0.630000 ;
      RECT 682.795000 0.000000 684.045000 0.630000 ;
      RECT 681.120000 0.000000 682.375000 0.630000 ;
      RECT 679.450000 0.000000 680.700000 0.630000 ;
      RECT 677.775000 0.000000 679.030000 0.630000 ;
      RECT 676.100000 0.000000 677.355000 0.630000 ;
      RECT 674.430000 0.000000 675.680000 0.630000 ;
      RECT 672.755000 0.000000 674.010000 0.630000 ;
      RECT 671.085000 0.000000 672.335000 0.630000 ;
      RECT 669.410000 0.000000 670.665000 0.630000 ;
      RECT 667.735000 0.000000 668.990000 0.630000 ;
      RECT 666.065000 0.000000 667.315000 0.630000 ;
      RECT 664.390000 0.000000 665.645000 0.630000 ;
      RECT 662.720000 0.000000 663.970000 0.630000 ;
      RECT 661.045000 0.000000 662.300000 0.630000 ;
      RECT 659.370000 0.000000 660.625000 0.630000 ;
      RECT 657.700000 0.000000 658.950000 0.630000 ;
      RECT 656.025000 0.000000 657.280000 0.630000 ;
      RECT 654.355000 0.000000 655.605000 0.630000 ;
      RECT 652.680000 0.000000 653.935000 0.630000 ;
      RECT 651.005000 0.000000 652.260000 0.630000 ;
      RECT 649.335000 0.000000 650.585000 0.630000 ;
      RECT 647.660000 0.000000 648.915000 0.630000 ;
      RECT 645.990000 0.000000 647.240000 0.630000 ;
      RECT 644.315000 0.000000 645.570000 0.630000 ;
      RECT 642.640000 0.000000 643.895000 0.630000 ;
      RECT 640.970000 0.000000 642.220000 0.630000 ;
      RECT 639.295000 0.000000 640.550000 0.630000 ;
      RECT 637.625000 0.000000 638.875000 0.630000 ;
      RECT 635.950000 0.000000 637.205000 0.630000 ;
      RECT 634.275000 0.000000 635.530000 0.630000 ;
      RECT 632.605000 0.000000 633.855000 0.630000 ;
      RECT 630.930000 0.000000 632.185000 0.630000 ;
      RECT 629.260000 0.000000 630.510000 0.630000 ;
      RECT 627.585000 0.000000 628.840000 0.630000 ;
      RECT 625.910000 0.000000 627.165000 0.630000 ;
      RECT 624.240000 0.000000 625.490000 0.630000 ;
      RECT 622.565000 0.000000 623.820000 0.630000 ;
      RECT 620.895000 0.000000 622.145000 0.630000 ;
      RECT 619.220000 0.000000 620.475000 0.630000 ;
      RECT 617.545000 0.000000 618.800000 0.630000 ;
      RECT 615.875000 0.000000 617.125000 0.630000 ;
      RECT 614.200000 0.000000 615.455000 0.630000 ;
      RECT 612.530000 0.000000 613.780000 0.630000 ;
      RECT 610.855000 0.000000 612.110000 0.630000 ;
      RECT 609.180000 0.000000 610.435000 0.630000 ;
      RECT 607.510000 0.000000 608.760000 0.630000 ;
      RECT 605.835000 0.000000 607.090000 0.630000 ;
      RECT 604.165000 0.000000 605.415000 0.630000 ;
      RECT 602.490000 0.000000 603.745000 0.630000 ;
      RECT 600.815000 0.000000 602.070000 0.630000 ;
      RECT 599.145000 0.000000 600.395000 0.630000 ;
      RECT 597.470000 0.000000 598.725000 0.630000 ;
      RECT 595.800000 0.000000 597.050000 0.630000 ;
      RECT 594.125000 0.000000 595.380000 0.630000 ;
      RECT 592.450000 0.000000 593.705000 0.630000 ;
      RECT 590.780000 0.000000 592.030000 0.630000 ;
      RECT 589.105000 0.000000 590.360000 0.630000 ;
      RECT 587.435000 0.000000 588.685000 0.630000 ;
      RECT 585.760000 0.000000 587.015000 0.630000 ;
      RECT 584.085000 0.000000 585.340000 0.630000 ;
      RECT 582.415000 0.000000 583.665000 0.630000 ;
      RECT 580.740000 0.000000 581.995000 0.630000 ;
      RECT 579.070000 0.000000 580.320000 0.630000 ;
      RECT 577.395000 0.000000 578.650000 0.630000 ;
      RECT 575.720000 0.000000 576.975000 0.630000 ;
      RECT 574.050000 0.000000 575.300000 0.630000 ;
      RECT 572.375000 0.000000 573.630000 0.630000 ;
      RECT 570.705000 0.000000 571.955000 0.630000 ;
      RECT 569.030000 0.000000 570.285000 0.630000 ;
      RECT 567.355000 0.000000 568.610000 0.630000 ;
      RECT 565.685000 0.000000 566.935000 0.630000 ;
      RECT 564.010000 0.000000 565.265000 0.630000 ;
      RECT 562.340000 0.000000 563.590000 0.630000 ;
      RECT 560.665000 0.000000 561.920000 0.630000 ;
      RECT 558.990000 0.000000 560.245000 0.630000 ;
      RECT 557.320000 0.000000 558.570000 0.630000 ;
      RECT 555.645000 0.000000 556.900000 0.630000 ;
      RECT 553.975000 0.000000 555.225000 0.630000 ;
      RECT 552.300000 0.000000 553.555000 0.630000 ;
      RECT 550.625000 0.000000 551.880000 0.630000 ;
      RECT 548.955000 0.000000 550.205000 0.630000 ;
      RECT 547.280000 0.000000 548.535000 0.630000 ;
      RECT 545.610000 0.000000 546.860000 0.630000 ;
      RECT 543.935000 0.000000 545.190000 0.630000 ;
      RECT 542.260000 0.000000 543.515000 0.630000 ;
      RECT 540.590000 0.000000 541.840000 0.630000 ;
      RECT 538.915000 0.000000 540.170000 0.630000 ;
      RECT 537.245000 0.000000 538.495000 0.630000 ;
      RECT 535.570000 0.000000 536.825000 0.630000 ;
      RECT 533.895000 0.000000 535.150000 0.630000 ;
      RECT 532.225000 0.000000 533.475000 0.630000 ;
      RECT 530.550000 0.000000 531.805000 0.630000 ;
      RECT 528.880000 0.000000 530.130000 0.630000 ;
      RECT 527.205000 0.000000 528.460000 0.630000 ;
      RECT 525.530000 0.000000 526.785000 0.630000 ;
      RECT 523.860000 0.000000 525.110000 0.630000 ;
      RECT 522.185000 0.000000 523.440000 0.630000 ;
      RECT 520.515000 0.000000 521.765000 0.630000 ;
      RECT 518.840000 0.000000 520.095000 0.630000 ;
      RECT 517.165000 0.000000 518.420000 0.630000 ;
      RECT 515.495000 0.000000 516.745000 0.630000 ;
      RECT 513.820000 0.000000 515.075000 0.630000 ;
      RECT 512.150000 0.000000 513.400000 0.630000 ;
      RECT 510.475000 0.000000 511.730000 0.630000 ;
      RECT 508.800000 0.000000 510.055000 0.630000 ;
      RECT 507.130000 0.000000 508.380000 0.630000 ;
      RECT 505.455000 0.000000 506.710000 0.630000 ;
      RECT 503.785000 0.000000 505.035000 0.630000 ;
      RECT 502.110000 0.000000 503.365000 0.630000 ;
      RECT 500.435000 0.000000 501.690000 0.630000 ;
      RECT 498.765000 0.000000 500.015000 0.630000 ;
      RECT 497.090000 0.000000 498.345000 0.630000 ;
      RECT 495.420000 0.000000 496.670000 0.630000 ;
      RECT 493.745000 0.000000 495.000000 0.630000 ;
      RECT 492.070000 0.000000 493.325000 0.630000 ;
      RECT 490.400000 0.000000 491.650000 0.630000 ;
      RECT 488.725000 0.000000 489.980000 0.630000 ;
      RECT 487.055000 0.000000 488.305000 0.630000 ;
      RECT 485.380000 0.000000 486.635000 0.630000 ;
      RECT 483.705000 0.000000 484.960000 0.630000 ;
      RECT 482.035000 0.000000 483.285000 0.630000 ;
      RECT 480.360000 0.000000 481.615000 0.630000 ;
      RECT 478.690000 0.000000 479.940000 0.630000 ;
      RECT 477.015000 0.000000 478.270000 0.630000 ;
      RECT 475.340000 0.000000 476.595000 0.630000 ;
      RECT 473.670000 0.000000 474.920000 0.630000 ;
      RECT 471.995000 0.000000 473.250000 0.630000 ;
      RECT 470.325000 0.000000 471.575000 0.630000 ;
      RECT 468.650000 0.000000 469.905000 0.630000 ;
      RECT 466.975000 0.000000 468.230000 0.630000 ;
      RECT 465.305000 0.000000 466.555000 0.630000 ;
      RECT 463.630000 0.000000 464.885000 0.630000 ;
      RECT 461.960000 0.000000 463.210000 0.630000 ;
      RECT 460.285000 0.000000 461.540000 0.630000 ;
      RECT 458.610000 0.000000 459.865000 0.630000 ;
      RECT 456.940000 0.000000 458.190000 0.630000 ;
      RECT 455.265000 0.000000 456.520000 0.630000 ;
      RECT 453.595000 0.000000 454.845000 0.630000 ;
      RECT 451.920000 0.000000 453.175000 0.630000 ;
      RECT 450.245000 0.000000 451.500000 0.630000 ;
      RECT 448.575000 0.000000 449.825000 0.630000 ;
      RECT 446.900000 0.000000 448.155000 0.630000 ;
      RECT 445.230000 0.000000 446.480000 0.630000 ;
      RECT 443.555000 0.000000 444.810000 0.630000 ;
      RECT 441.880000 0.000000 443.135000 0.630000 ;
      RECT 440.210000 0.000000 441.460000 0.630000 ;
      RECT 438.535000 0.000000 439.790000 0.630000 ;
      RECT 436.865000 0.000000 438.115000 0.630000 ;
      RECT 435.190000 0.000000 436.445000 0.630000 ;
      RECT 433.515000 0.000000 434.770000 0.630000 ;
      RECT 431.845000 0.000000 433.095000 0.630000 ;
      RECT 430.170000 0.000000 431.425000 0.630000 ;
      RECT 428.500000 0.000000 429.750000 0.630000 ;
      RECT 426.825000 0.000000 428.080000 0.630000 ;
      RECT 425.150000 0.000000 426.405000 0.630000 ;
      RECT 423.480000 0.000000 424.730000 0.630000 ;
      RECT 421.805000 0.000000 423.060000 0.630000 ;
      RECT 420.135000 0.000000 421.385000 0.630000 ;
      RECT 418.460000 0.000000 419.715000 0.630000 ;
      RECT 416.785000 0.000000 418.040000 0.630000 ;
      RECT 415.115000 0.000000 416.365000 0.630000 ;
      RECT 413.440000 0.000000 414.695000 0.630000 ;
      RECT 411.770000 0.000000 413.020000 0.630000 ;
      RECT 410.095000 0.000000 411.350000 0.630000 ;
      RECT 408.420000 0.000000 409.675000 0.630000 ;
      RECT 406.750000 0.000000 408.000000 0.630000 ;
      RECT 405.075000 0.000000 406.330000 0.630000 ;
      RECT 403.405000 0.000000 404.655000 0.630000 ;
      RECT 401.730000 0.000000 402.985000 0.630000 ;
      RECT 400.055000 0.000000 401.310000 0.630000 ;
      RECT 398.385000 0.000000 399.635000 0.630000 ;
      RECT 396.710000 0.000000 397.965000 0.630000 ;
      RECT 395.040000 0.000000 396.290000 0.630000 ;
      RECT 393.365000 0.000000 394.620000 0.630000 ;
      RECT 391.690000 0.000000 392.945000 0.630000 ;
      RECT 390.020000 0.000000 391.270000 0.630000 ;
      RECT 388.345000 0.000000 389.600000 0.630000 ;
      RECT 386.675000 0.000000 387.925000 0.630000 ;
      RECT 385.000000 0.000000 386.255000 0.630000 ;
      RECT 383.325000 0.000000 384.580000 0.630000 ;
      RECT 381.655000 0.000000 382.905000 0.630000 ;
      RECT 379.980000 0.000000 381.235000 0.630000 ;
      RECT 378.310000 0.000000 379.560000 0.630000 ;
      RECT 376.635000 0.000000 377.890000 0.630000 ;
      RECT 374.960000 0.000000 376.215000 0.630000 ;
      RECT 373.290000 0.000000 374.540000 0.630000 ;
      RECT 371.615000 0.000000 372.870000 0.630000 ;
      RECT 369.945000 0.000000 371.195000 0.630000 ;
      RECT 368.270000 0.000000 369.525000 0.630000 ;
      RECT 366.595000 0.000000 367.850000 0.630000 ;
      RECT 364.925000 0.000000 366.175000 0.630000 ;
      RECT 363.250000 0.000000 364.505000 0.630000 ;
      RECT 361.580000 0.000000 362.830000 0.630000 ;
      RECT 359.905000 0.000000 361.160000 0.630000 ;
      RECT 358.230000 0.000000 359.485000 0.630000 ;
      RECT 356.560000 0.000000 357.810000 0.630000 ;
      RECT 354.885000 0.000000 356.140000 0.630000 ;
      RECT 353.215000 0.000000 354.465000 0.630000 ;
      RECT 351.540000 0.000000 352.795000 0.630000 ;
      RECT 349.865000 0.000000 351.120000 0.630000 ;
      RECT 348.195000 0.000000 349.445000 0.630000 ;
      RECT 346.520000 0.000000 347.775000 0.630000 ;
      RECT 344.850000 0.000000 346.100000 0.630000 ;
      RECT 343.175000 0.000000 344.430000 0.630000 ;
      RECT 341.500000 0.000000 342.755000 0.630000 ;
      RECT 339.830000 0.000000 341.080000 0.630000 ;
      RECT 338.155000 0.000000 339.410000 0.630000 ;
      RECT 336.485000 0.000000 337.735000 0.630000 ;
      RECT 334.810000 0.000000 336.065000 0.630000 ;
      RECT 333.135000 0.000000 334.390000 0.630000 ;
      RECT 331.465000 0.000000 332.715000 0.630000 ;
      RECT 329.790000 0.000000 331.045000 0.630000 ;
      RECT 328.120000 0.000000 329.370000 0.630000 ;
      RECT 326.445000 0.000000 327.700000 0.630000 ;
      RECT 324.770000 0.000000 326.025000 0.630000 ;
      RECT 323.100000 0.000000 324.350000 0.630000 ;
      RECT 321.425000 0.000000 322.680000 0.630000 ;
      RECT 319.755000 0.000000 321.005000 0.630000 ;
      RECT 318.080000 0.000000 319.335000 0.630000 ;
      RECT 316.405000 0.000000 317.660000 0.630000 ;
      RECT 314.735000 0.000000 315.985000 0.630000 ;
      RECT 313.060000 0.000000 314.315000 0.630000 ;
      RECT 311.390000 0.000000 312.640000 0.630000 ;
      RECT 309.715000 0.000000 310.970000 0.630000 ;
      RECT 308.040000 0.000000 309.295000 0.630000 ;
      RECT 306.370000 0.000000 307.620000 0.630000 ;
      RECT 304.695000 0.000000 305.950000 0.630000 ;
      RECT 303.025000 0.000000 304.275000 0.630000 ;
      RECT 301.350000 0.000000 302.605000 0.630000 ;
      RECT 299.675000 0.000000 300.930000 0.630000 ;
      RECT 298.005000 0.000000 299.255000 0.630000 ;
      RECT 296.330000 0.000000 297.585000 0.630000 ;
      RECT 294.660000 0.000000 295.910000 0.630000 ;
      RECT 292.985000 0.000000 294.240000 0.630000 ;
      RECT 291.310000 0.000000 292.565000 0.630000 ;
      RECT 289.640000 0.000000 290.890000 0.630000 ;
      RECT 287.965000 0.000000 289.220000 0.630000 ;
      RECT 286.295000 0.000000 287.545000 0.630000 ;
      RECT 284.620000 0.000000 285.875000 0.630000 ;
      RECT 282.945000 0.000000 284.200000 0.630000 ;
      RECT 281.275000 0.000000 282.525000 0.630000 ;
      RECT 279.600000 0.000000 280.855000 0.630000 ;
      RECT 277.930000 0.000000 279.180000 0.630000 ;
      RECT 276.255000 0.000000 277.510000 0.630000 ;
      RECT 274.580000 0.000000 275.835000 0.630000 ;
      RECT 272.910000 0.000000 274.160000 0.630000 ;
      RECT 271.235000 0.000000 272.490000 0.630000 ;
      RECT 269.565000 0.000000 270.815000 0.630000 ;
      RECT 267.890000 0.000000 269.145000 0.630000 ;
      RECT 266.215000 0.000000 267.470000 0.630000 ;
      RECT 264.545000 0.000000 265.795000 0.630000 ;
      RECT 262.870000 0.000000 264.125000 0.630000 ;
      RECT 261.200000 0.000000 262.450000 0.630000 ;
      RECT 259.525000 0.000000 260.780000 0.630000 ;
      RECT 257.850000 0.000000 259.105000 0.630000 ;
      RECT 256.180000 0.000000 257.430000 0.630000 ;
      RECT 254.505000 0.000000 255.760000 0.630000 ;
      RECT 252.835000 0.000000 254.085000 0.630000 ;
      RECT 251.160000 0.000000 252.415000 0.630000 ;
      RECT 249.485000 0.000000 250.740000 0.630000 ;
      RECT 247.815000 0.000000 249.065000 0.630000 ;
      RECT 246.140000 0.000000 247.395000 0.630000 ;
      RECT 244.470000 0.000000 245.720000 0.630000 ;
      RECT 242.795000 0.000000 244.050000 0.630000 ;
      RECT 241.120000 0.000000 242.375000 0.630000 ;
      RECT 239.450000 0.000000 240.700000 0.630000 ;
      RECT 237.775000 0.000000 239.030000 0.630000 ;
      RECT 236.105000 0.000000 237.355000 0.630000 ;
      RECT 234.430000 0.000000 235.685000 0.630000 ;
      RECT 232.755000 0.000000 234.010000 0.630000 ;
      RECT 231.085000 0.000000 232.335000 0.630000 ;
      RECT 229.410000 0.000000 230.665000 0.630000 ;
      RECT 227.740000 0.000000 228.990000 0.630000 ;
      RECT 226.065000 0.000000 227.320000 0.630000 ;
      RECT 224.390000 0.000000 225.645000 0.630000 ;
      RECT 222.720000 0.000000 223.970000 0.630000 ;
      RECT 221.045000 0.000000 222.300000 0.630000 ;
      RECT 219.375000 0.000000 220.625000 0.630000 ;
      RECT 217.700000 0.000000 218.955000 0.630000 ;
      RECT 216.025000 0.000000 217.280000 0.630000 ;
      RECT 214.355000 0.000000 215.605000 0.630000 ;
      RECT 212.680000 0.000000 213.935000 0.630000 ;
      RECT 211.010000 0.000000 212.260000 0.630000 ;
      RECT 209.335000 0.000000 210.590000 0.630000 ;
      RECT 207.660000 0.000000 208.915000 0.630000 ;
      RECT 205.990000 0.000000 207.240000 0.630000 ;
      RECT 204.315000 0.000000 205.570000 0.630000 ;
      RECT 202.645000 0.000000 203.895000 0.630000 ;
      RECT 200.970000 0.000000 202.225000 0.630000 ;
      RECT 199.295000 0.000000 200.550000 0.630000 ;
      RECT 197.625000 0.000000 198.875000 0.630000 ;
      RECT 195.950000 0.000000 197.205000 0.630000 ;
      RECT 194.280000 0.000000 195.530000 0.630000 ;
      RECT 192.605000 0.000000 193.860000 0.630000 ;
      RECT 190.930000 0.000000 192.185000 0.630000 ;
      RECT 189.260000 0.000000 190.510000 0.630000 ;
      RECT 187.585000 0.000000 188.840000 0.630000 ;
      RECT 185.915000 0.000000 187.165000 0.630000 ;
      RECT 184.240000 0.000000 185.495000 0.630000 ;
      RECT 182.565000 0.000000 183.820000 0.630000 ;
      RECT 180.895000 0.000000 182.145000 0.630000 ;
      RECT 179.220000 0.000000 180.475000 0.630000 ;
      RECT 177.550000 0.000000 178.800000 0.630000 ;
      RECT 175.875000 0.000000 177.130000 0.630000 ;
      RECT 174.200000 0.000000 175.455000 0.630000 ;
      RECT 172.530000 0.000000 173.780000 0.630000 ;
      RECT 170.855000 0.000000 172.110000 0.630000 ;
      RECT 169.185000 0.000000 170.435000 0.630000 ;
      RECT 167.510000 0.000000 168.765000 0.630000 ;
      RECT 165.835000 0.000000 167.090000 0.630000 ;
      RECT 164.165000 0.000000 165.415000 0.630000 ;
      RECT 162.490000 0.000000 163.745000 0.630000 ;
      RECT 160.820000 0.000000 162.070000 0.630000 ;
      RECT 159.145000 0.000000 160.400000 0.630000 ;
      RECT 157.470000 0.000000 158.725000 0.630000 ;
      RECT 155.800000 0.000000 157.050000 0.630000 ;
      RECT 154.125000 0.000000 155.380000 0.630000 ;
      RECT 152.455000 0.000000 153.705000 0.630000 ;
      RECT 150.780000 0.000000 152.035000 0.630000 ;
      RECT 149.105000 0.000000 150.360000 0.630000 ;
      RECT 147.435000 0.000000 148.685000 0.630000 ;
      RECT 145.760000 0.000000 147.015000 0.630000 ;
      RECT 144.090000 0.000000 145.340000 0.630000 ;
      RECT 142.415000 0.000000 143.670000 0.630000 ;
      RECT 140.740000 0.000000 141.995000 0.630000 ;
      RECT 139.070000 0.000000 140.320000 0.630000 ;
      RECT 137.395000 0.000000 138.650000 0.630000 ;
      RECT 135.725000 0.000000 136.975000 0.630000 ;
      RECT 134.050000 0.000000 135.305000 0.630000 ;
      RECT 132.375000 0.000000 133.630000 0.630000 ;
      RECT 130.705000 0.000000 131.955000 0.630000 ;
      RECT 129.030000 0.000000 130.285000 0.630000 ;
      RECT 127.360000 0.000000 128.610000 0.630000 ;
      RECT 125.685000 0.000000 126.940000 0.630000 ;
      RECT 124.010000 0.000000 125.265000 0.630000 ;
      RECT 122.340000 0.000000 123.590000 0.630000 ;
      RECT 120.665000 0.000000 121.920000 0.630000 ;
      RECT 118.995000 0.000000 120.245000 0.630000 ;
      RECT 117.320000 0.000000 118.575000 0.630000 ;
      RECT 115.645000 0.000000 116.900000 0.630000 ;
      RECT 113.975000 0.000000 115.225000 0.630000 ;
      RECT 112.300000 0.000000 113.555000 0.630000 ;
      RECT 110.630000 0.000000 111.880000 0.630000 ;
      RECT 108.955000 0.000000 110.210000 0.630000 ;
      RECT 107.280000 0.000000 108.535000 0.630000 ;
      RECT 105.610000 0.000000 106.860000 0.630000 ;
      RECT 103.935000 0.000000 105.190000 0.630000 ;
      RECT 102.265000 0.000000 103.515000 0.630000 ;
      RECT 100.590000 0.000000 101.845000 0.630000 ;
      RECT 98.915000 0.000000 100.170000 0.630000 ;
      RECT 97.245000 0.000000 98.495000 0.630000 ;
      RECT 95.570000 0.000000 96.825000 0.630000 ;
      RECT 93.900000 0.000000 95.150000 0.630000 ;
      RECT 92.225000 0.000000 93.480000 0.630000 ;
      RECT 90.550000 0.000000 91.805000 0.630000 ;
      RECT 88.880000 0.000000 90.130000 0.630000 ;
      RECT 87.205000 0.000000 88.460000 0.630000 ;
      RECT 85.535000 0.000000 86.785000 0.630000 ;
      RECT 83.860000 0.000000 85.115000 0.630000 ;
      RECT 82.185000 0.000000 83.440000 0.630000 ;
      RECT 80.515000 0.000000 81.765000 0.630000 ;
      RECT 78.840000 0.000000 80.095000 0.630000 ;
      RECT 77.170000 0.000000 78.420000 0.630000 ;
      RECT 75.495000 0.000000 76.750000 0.630000 ;
      RECT 73.820000 0.000000 75.075000 0.630000 ;
      RECT 72.150000 0.000000 73.400000 0.630000 ;
      RECT 70.475000 0.000000 71.730000 0.630000 ;
      RECT 68.805000 0.000000 70.055000 0.630000 ;
      RECT 67.130000 0.000000 68.385000 0.630000 ;
      RECT 65.455000 0.000000 66.710000 0.630000 ;
      RECT 63.785000 0.000000 65.035000 0.630000 ;
      RECT 62.110000 0.000000 63.365000 0.630000 ;
      RECT 60.440000 0.000000 61.690000 0.630000 ;
      RECT 58.765000 0.000000 60.020000 0.630000 ;
      RECT 57.090000 0.000000 58.345000 0.630000 ;
      RECT 55.420000 0.000000 56.670000 0.630000 ;
      RECT 53.745000 0.000000 55.000000 0.630000 ;
      RECT 52.075000 0.000000 53.325000 0.630000 ;
      RECT 50.400000 0.000000 51.655000 0.630000 ;
      RECT 48.725000 0.000000 49.980000 0.630000 ;
      RECT 47.055000 0.000000 48.305000 0.630000 ;
      RECT 45.380000 0.000000 46.635000 0.630000 ;
      RECT 43.710000 0.000000 44.960000 0.630000 ;
      RECT 42.035000 0.000000 43.290000 0.630000 ;
      RECT 40.360000 0.000000 41.615000 0.630000 ;
      RECT 38.690000 0.000000 39.940000 0.630000 ;
      RECT 37.015000 0.000000 38.270000 0.630000 ;
      RECT 35.345000 0.000000 36.595000 0.630000 ;
      RECT 33.670000 0.000000 34.925000 0.630000 ;
      RECT 31.995000 0.000000 33.250000 0.630000 ;
      RECT 30.325000 0.000000 31.575000 0.630000 ;
      RECT 28.650000 0.000000 29.905000 0.630000 ;
      RECT 26.980000 0.000000 28.230000 0.630000 ;
      RECT 25.305000 0.000000 26.560000 0.630000 ;
      RECT 23.630000 0.000000 24.885000 0.630000 ;
      RECT 21.960000 0.000000 23.210000 0.630000 ;
      RECT 20.285000 0.000000 21.540000 0.630000 ;
      RECT 18.615000 0.000000 19.865000 0.630000 ;
      RECT 16.940000 0.000000 18.195000 0.630000 ;
      RECT 15.265000 0.000000 16.520000 0.630000 ;
      RECT 13.595000 0.000000 14.845000 0.630000 ;
      RECT 11.920000 0.000000 13.175000 0.630000 ;
      RECT 10.250000 0.000000 11.500000 0.630000 ;
      RECT 8.575000 0.000000 9.830000 0.630000 ;
      RECT 6.900000 0.000000 8.155000 0.630000 ;
      RECT 5.230000 0.000000 6.480000 0.630000 ;
      RECT 3.555000 0.000000 4.810000 0.630000 ;
      RECT 1.885000 0.000000 3.135000 0.630000 ;
      RECT 0.900000 0.000000 1.465000 0.630000 ;
      RECT 0.000000 0.000000 0.480000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 811.140000 818.340000 814.640000 ;
      RECT 1.100000 810.530000 818.340000 811.140000 ;
      RECT 1.100000 810.240000 817.240000 810.530000 ;
      RECT 0.000000 809.630000 817.240000 810.240000 ;
      RECT 0.000000 796.550000 818.340000 809.630000 ;
      RECT 0.000000 795.650000 817.240000 796.550000 ;
      RECT 0.000000 795.210000 818.340000 795.650000 ;
      RECT 1.100000 794.310000 818.340000 795.210000 ;
      RECT 0.000000 778.040000 818.340000 794.310000 ;
      RECT 0.000000 777.140000 817.240000 778.040000 ;
      RECT 0.000000 775.340000 818.340000 777.140000 ;
      RECT 1.100000 774.440000 818.340000 775.340000 ;
      RECT 0.000000 759.525000 818.340000 774.440000 ;
      RECT 0.000000 758.625000 817.240000 759.525000 ;
      RECT 0.000000 755.470000 818.340000 758.625000 ;
      RECT 1.100000 754.570000 818.340000 755.470000 ;
      RECT 0.000000 741.010000 818.340000 754.570000 ;
      RECT 0.000000 740.110000 817.240000 741.010000 ;
      RECT 0.000000 735.605000 818.340000 740.110000 ;
      RECT 1.100000 734.705000 818.340000 735.605000 ;
      RECT 0.000000 722.495000 818.340000 734.705000 ;
      RECT 0.000000 721.595000 817.240000 722.495000 ;
      RECT 0.000000 715.735000 818.340000 721.595000 ;
      RECT 1.100000 714.835000 818.340000 715.735000 ;
      RECT 0.000000 703.980000 818.340000 714.835000 ;
      RECT 0.000000 703.080000 817.240000 703.980000 ;
      RECT 0.000000 695.865000 818.340000 703.080000 ;
      RECT 1.100000 694.965000 818.340000 695.865000 ;
      RECT 0.000000 685.470000 818.340000 694.965000 ;
      RECT 0.000000 684.570000 817.240000 685.470000 ;
      RECT 0.000000 675.995000 818.340000 684.570000 ;
      RECT 1.100000 675.095000 818.340000 675.995000 ;
      RECT 0.000000 666.955000 818.340000 675.095000 ;
      RECT 0.000000 666.055000 817.240000 666.955000 ;
      RECT 0.000000 656.125000 818.340000 666.055000 ;
      RECT 1.100000 655.225000 818.340000 656.125000 ;
      RECT 0.000000 648.440000 818.340000 655.225000 ;
      RECT 0.000000 647.540000 817.240000 648.440000 ;
      RECT 0.000000 636.260000 818.340000 647.540000 ;
      RECT 1.100000 635.360000 818.340000 636.260000 ;
      RECT 0.000000 629.925000 818.340000 635.360000 ;
      RECT 0.000000 629.025000 817.240000 629.925000 ;
      RECT 0.000000 616.390000 818.340000 629.025000 ;
      RECT 1.100000 615.490000 818.340000 616.390000 ;
      RECT 0.000000 611.410000 818.340000 615.490000 ;
      RECT 0.000000 610.510000 817.240000 611.410000 ;
      RECT 0.000000 596.520000 818.340000 610.510000 ;
      RECT 1.100000 595.620000 818.340000 596.520000 ;
      RECT 0.000000 592.900000 818.340000 595.620000 ;
      RECT 0.000000 592.000000 817.240000 592.900000 ;
      RECT 0.000000 576.650000 818.340000 592.000000 ;
      RECT 1.100000 575.750000 818.340000 576.650000 ;
      RECT 0.000000 574.385000 818.340000 575.750000 ;
      RECT 0.000000 573.485000 817.240000 574.385000 ;
      RECT 0.000000 556.780000 818.340000 573.485000 ;
      RECT 1.100000 555.880000 818.340000 556.780000 ;
      RECT 0.000000 555.870000 818.340000 555.880000 ;
      RECT 0.000000 554.970000 817.240000 555.870000 ;
      RECT 0.000000 537.355000 818.340000 554.970000 ;
      RECT 0.000000 536.915000 817.240000 537.355000 ;
      RECT 1.100000 536.455000 817.240000 536.915000 ;
      RECT 1.100000 536.015000 818.340000 536.455000 ;
      RECT 0.000000 518.840000 818.340000 536.015000 ;
      RECT 0.000000 517.940000 817.240000 518.840000 ;
      RECT 0.000000 517.045000 818.340000 517.940000 ;
      RECT 1.100000 516.145000 818.340000 517.045000 ;
      RECT 0.000000 500.330000 818.340000 516.145000 ;
      RECT 0.000000 499.430000 817.240000 500.330000 ;
      RECT 0.000000 497.175000 818.340000 499.430000 ;
      RECT 1.100000 496.275000 818.340000 497.175000 ;
      RECT 0.000000 481.815000 818.340000 496.275000 ;
      RECT 0.000000 480.915000 817.240000 481.815000 ;
      RECT 0.000000 477.305000 818.340000 480.915000 ;
      RECT 1.100000 476.405000 818.340000 477.305000 ;
      RECT 0.000000 463.300000 818.340000 476.405000 ;
      RECT 0.000000 462.400000 817.240000 463.300000 ;
      RECT 0.000000 457.435000 818.340000 462.400000 ;
      RECT 1.100000 456.535000 818.340000 457.435000 ;
      RECT 0.000000 444.785000 818.340000 456.535000 ;
      RECT 0.000000 443.885000 817.240000 444.785000 ;
      RECT 0.000000 437.570000 818.340000 443.885000 ;
      RECT 1.100000 436.670000 818.340000 437.570000 ;
      RECT 0.000000 426.270000 818.340000 436.670000 ;
      RECT 0.000000 425.370000 817.240000 426.270000 ;
      RECT 0.000000 417.700000 818.340000 425.370000 ;
      RECT 1.100000 416.800000 818.340000 417.700000 ;
      RECT 0.000000 407.760000 818.340000 416.800000 ;
      RECT 0.000000 406.860000 817.240000 407.760000 ;
      RECT 0.000000 397.830000 818.340000 406.860000 ;
      RECT 1.100000 396.930000 818.340000 397.830000 ;
      RECT 0.000000 389.245000 818.340000 396.930000 ;
      RECT 0.000000 388.345000 817.240000 389.245000 ;
      RECT 0.000000 377.960000 818.340000 388.345000 ;
      RECT 1.100000 377.060000 818.340000 377.960000 ;
      RECT 0.000000 370.730000 818.340000 377.060000 ;
      RECT 0.000000 369.830000 817.240000 370.730000 ;
      RECT 0.000000 358.090000 818.340000 369.830000 ;
      RECT 1.100000 357.190000 818.340000 358.090000 ;
      RECT 0.000000 352.215000 818.340000 357.190000 ;
      RECT 0.000000 351.315000 817.240000 352.215000 ;
      RECT 0.000000 338.225000 818.340000 351.315000 ;
      RECT 1.100000 337.325000 818.340000 338.225000 ;
      RECT 0.000000 333.700000 818.340000 337.325000 ;
      RECT 0.000000 332.800000 817.240000 333.700000 ;
      RECT 0.000000 318.355000 818.340000 332.800000 ;
      RECT 1.100000 317.455000 818.340000 318.355000 ;
      RECT 0.000000 315.190000 818.340000 317.455000 ;
      RECT 0.000000 314.290000 817.240000 315.190000 ;
      RECT 0.000000 298.485000 818.340000 314.290000 ;
      RECT 1.100000 297.585000 818.340000 298.485000 ;
      RECT 0.000000 296.675000 818.340000 297.585000 ;
      RECT 0.000000 295.775000 817.240000 296.675000 ;
      RECT 0.000000 278.615000 818.340000 295.775000 ;
      RECT 1.100000 278.160000 818.340000 278.615000 ;
      RECT 1.100000 277.715000 817.240000 278.160000 ;
      RECT 0.000000 277.260000 817.240000 277.715000 ;
      RECT 0.000000 259.645000 818.340000 277.260000 ;
      RECT 0.000000 258.745000 817.240000 259.645000 ;
      RECT 1.100000 257.845000 818.340000 258.745000 ;
      RECT 0.000000 241.130000 818.340000 257.845000 ;
      RECT 0.000000 240.230000 817.240000 241.130000 ;
      RECT 0.000000 238.880000 818.340000 240.230000 ;
      RECT 1.100000 237.980000 818.340000 238.880000 ;
      RECT 0.000000 222.620000 818.340000 237.980000 ;
      RECT 0.000000 221.720000 817.240000 222.620000 ;
      RECT 0.000000 219.010000 818.340000 221.720000 ;
      RECT 1.100000 218.110000 818.340000 219.010000 ;
      RECT 0.000000 204.105000 818.340000 218.110000 ;
      RECT 0.000000 203.205000 817.240000 204.105000 ;
      RECT 0.000000 199.140000 818.340000 203.205000 ;
      RECT 1.100000 198.240000 818.340000 199.140000 ;
      RECT 0.000000 185.590000 818.340000 198.240000 ;
      RECT 0.000000 184.690000 817.240000 185.590000 ;
      RECT 0.000000 179.270000 818.340000 184.690000 ;
      RECT 1.100000 178.370000 818.340000 179.270000 ;
      RECT 0.000000 167.075000 818.340000 178.370000 ;
      RECT 0.000000 166.175000 817.240000 167.075000 ;
      RECT 0.000000 159.400000 818.340000 166.175000 ;
      RECT 1.100000 158.500000 818.340000 159.400000 ;
      RECT 0.000000 148.560000 818.340000 158.500000 ;
      RECT 0.000000 147.660000 817.240000 148.560000 ;
      RECT 0.000000 139.535000 818.340000 147.660000 ;
      RECT 1.100000 138.635000 818.340000 139.535000 ;
      RECT 0.000000 130.050000 818.340000 138.635000 ;
      RECT 0.000000 129.150000 817.240000 130.050000 ;
      RECT 0.000000 119.665000 818.340000 129.150000 ;
      RECT 1.100000 118.765000 818.340000 119.665000 ;
      RECT 0.000000 111.535000 818.340000 118.765000 ;
      RECT 0.000000 110.635000 817.240000 111.535000 ;
      RECT 0.000000 99.795000 818.340000 110.635000 ;
      RECT 1.100000 98.895000 818.340000 99.795000 ;
      RECT 0.000000 93.020000 818.340000 98.895000 ;
      RECT 0.000000 92.120000 817.240000 93.020000 ;
      RECT 0.000000 79.925000 818.340000 92.120000 ;
      RECT 1.100000 79.025000 818.340000 79.925000 ;
      RECT 0.000000 74.505000 818.340000 79.025000 ;
      RECT 0.000000 73.605000 817.240000 74.505000 ;
      RECT 0.000000 60.055000 818.340000 73.605000 ;
      RECT 1.100000 59.155000 818.340000 60.055000 ;
      RECT 0.000000 55.990000 818.340000 59.155000 ;
      RECT 0.000000 55.090000 817.240000 55.990000 ;
      RECT 0.000000 40.190000 818.340000 55.090000 ;
      RECT 1.100000 39.290000 818.340000 40.190000 ;
      RECT 0.000000 37.480000 818.340000 39.290000 ;
      RECT 0.000000 36.580000 817.240000 37.480000 ;
      RECT 0.000000 20.320000 818.340000 36.580000 ;
      RECT 1.100000 19.420000 818.340000 20.320000 ;
      RECT 0.000000 18.965000 818.340000 19.420000 ;
      RECT 0.000000 18.065000 817.240000 18.965000 ;
      RECT 0.000000 10.820000 818.340000 18.065000 ;
      RECT 1.100000 10.210000 818.340000 10.820000 ;
      RECT 1.100000 9.920000 817.240000 10.210000 ;
      RECT 0.000000 9.310000 817.240000 9.920000 ;
      RECT 0.000000 0.000000 818.340000 9.310000 ;
    LAYER met4 ;
      RECT 0.000000 814.340000 818.340000 814.640000 ;
      RECT 2.860000 807.340000 815.480000 814.340000 ;
      RECT 811.080000 7.300000 815.480000 807.340000 ;
      RECT 9.860000 7.300000 808.480000 807.340000 ;
      RECT 2.860000 7.300000 7.260000 807.340000 ;
      RECT 818.080000 0.300000 818.340000 814.340000 ;
      RECT 2.860000 0.300000 815.480000 7.300000 ;
      RECT 0.000000 0.300000 0.260000 814.340000 ;
      RECT 0.000000 0.000000 818.340000 0.300000 ;
  END
END user_proj_example

END LIBRARY
